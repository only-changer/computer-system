/* ACM Class System (I) 2017 Fall Homework 1 
 *
 * PART II: Correct the following program
 * 
 * GUIDE:
 *   1. Create a RTL project in Vivado
 *   2. Put this file into `Simulation Sources'
 *   3. Run Behavioral Simulation
 *   4. You can see the results in `Tcl console'
 *
 */

module testfault;
	reg[15:0] a,b;
	wire[15:0] answer;
	fault f(a,b,answer);
	initial begin
		a = 10;
		b = 20;
		
		#1;
		if(answer != 20) begin
			$display("Expected 20, got %d", answer);
			$fatal("Wrong Answer");
		end
		
		#1;
		
		a = 40;
		b = 30;
		
		#1;
		
		if(answer != 40) begin
			$display("Expected 40, got %d", answer);
			$fatal("Wrong Answer");
		end
		
		$display("Congratulations! You have passed this test.");
		$finish;
	end
endmodule

module fault(a,b,answer);
	input wire[15:0] a,b;
	output wire[15:0] answer;
	wire [15 : 0] c;
	wire [15 : 0] d;
	assign c[15] = (! a[15]) & b[15];
	assign d[15] = (! a[15]) | b[15];
	assign answer[15] = a[15] | b[15];
	
	assign answer[14] = ((c[15] ^ d[15]) & (a[14] | b[14])) | ((!(c[15] ^ d[15])) & c[15] & d[15] & b[14]) | ((!(c[15] ^ d[15])) & (!(c[15] & d[15])) & a[14]);
	assign c[14] = ((c[15] ^ d[15]) & (! a[14]) & b[14]) | ((!(c[15] ^ d[15])) & c[15] & d[15] & 1) | ((!(c[15] ^ d[15])) & (!(c[15] & d[15])) & 0);
	assign d[14] = ((c[15] ^ d[15]) & ((! a[14]) | b[14])) | ((!(c[15] ^ d[15])) & c[15] & d[15] & 1) | ((!(c[15] ^ d[15])) & (!(c[15] & d[15])) & 0);
	
	assign answer[13] = ((c[14] ^ d[14]) & (a[13] | b[13])) | ((!(c[14] ^ d[14])) & c[14] & d[14] & b[13]) | ((!(c[14] ^ d[14])) & (!(c[14] & d[14])) & a[13]);
    assign c[13] = ((c[14] ^ d[14]) & (! a[13]) & b[13]) | ((!(c[14] ^ d[14])) & c[14] & d[14] & 1) | ((!(c[14] ^ d[14])) & (!(c[14] & d[14])) & 0);
    assign d[13] = ((c[14] ^ d[14]) & ((! a[13]) | b[13])) | ((!(c[14] ^ d[14])) & c[14] & d[14] & 1) | ((!(c[14] ^ d[14])) & (!(c[14] & d[14])) & 0);
    
    assign answer[12] = ((c[13] ^ d[13]) & (a[12] | b[12])) | ((!(c[13] ^ d[13])) & c[13] & d[13] & b[12]) | ((!(c[13] ^ d[13])) & (!(c[13] & d[13])) & a[12]);
    assign c[12] = ((c[13] ^ d[13]) & (! a[12]) & b[12]) | ((!(c[13] ^ d[13])) & c[13] & d[13] & 1) | ((!(c[13] ^ d[13])) & (!(c[13] & d[13])) & 0);
    assign d[12] = ((c[13] ^ d[13]) & ((! a[12]) | b[12])) | ((!(c[13] ^ d[13])) & c[13] & d[13] & 1) | ((!(c[13] ^ d[13])) & (!(c[13] & d[13])) & 0);
    
    assign answer[11] = ((c[12] ^ d[12]) & (a[11] | b[11])) | ((!(c[12] ^ d[12])) & c[12] & d[12] & b[11]) | ((!(c[12] ^ d[12])) & (!(c[12] & d[12])) & a[11]);
    assign c[11] = ((c[12] ^ d[12]) & (! a[11]) & b[11]) | ((!(c[12] ^ d[12])) & c[12] & d[12] & 1) | ((!(c[12] ^ d[12])) & (!(c[12] & d[12])) & 0);
    assign d[11] = ((c[12] ^ d[12]) & ((! a[11]) | b[11])) | ((!(c[12] ^ d[12])) & c[12] & d[12] & 1) | ((!(c[12] ^ d[12])) & (!(c[12] & d[12])) & 0);
    
    assign answer[10] = ((c[11] ^ d[11]) & (a[10] | b[10])) | ((!(c[11] ^ d[11])) & c[11] & d[11] & b[10]) | ((!(c[11] ^ d[11])) & (!(c[11] & d[11])) & a[10]);
    assign c[10] = ((c[11] ^ d[11]) & (! a[10]) & b[10]) | ((!(c[11] ^ d[11])) & c[11] & d[11] & 1) | ((!(c[11] ^ d[11])) & (!(c[11] & d[11])) & 0);
    assign d[10] = ((c[11] ^ d[11]) & ((! a[10]) | b[10])) | ((!(c[11] ^ d[11])) & c[11] & d[11] & 1) | ((!(c[11] ^ d[11])) & (!(c[11] & d[11])) & 0);
    
    assign answer[9] = ((c[10] ^ d[10]) & (a[9] | b[9])) | ((!(c[10] ^ d[10])) & c[10] & d[10] & b[9]) | ((!(c[10] ^ d[10])) & (!(c[10] & d[10])) & a[9]);
    assign c[9] = ((c[10] ^ d[10]) & (! a[9]) & b[9]) | ((!(c[10] ^ d[10])) & c[10] & d[10] & 1) | ((!(c[10] ^ d[10])) & (!(c[10] & d[10])) & 0);
    assign d[9] = ((c[10] ^ d[10]) & ((! a[9]) | b[9])) | ((!(c[10] ^ d[10])) & c[10] & d[10] & 1) | ((!(c[10] ^ d[10])) & (!(c[10] & d[10])) & 0);
    
    assign answer[8] = ((c[9] ^ d[9]) & (a[8] | b[8])) | ((!(c[9] ^ d[9])) & c[9] & d[9] & b[8]) | ((!(c[9] ^ d[9])) & (!(c[9] & d[9])) & a[8]);
    assign c[8] = ((c[9] ^ d[9]) & (! a[8]) & b[8]) | ((!(c[9] ^ d[9])) & c[9] & d[9] & 1) | ((!(c[9] ^ d[9])) & (!(c[9] & d[9])) & 0);
    assign d[8] = ((c[9] ^ d[9]) & ((! a[8]) | b[8])) | ((!(c[9] ^ d[9])) & c[9] & d[9] & 1) | ((!(c[9] ^ d[9])) & (!(c[9] & d[9])) & 0);
    
    assign answer[7] = ((c[8] ^ d[8]) & (a[7] | b[7])) | ((!(c[8] ^ d[8])) & c[8] & d[8] & b[7]) | ((!(c[8] ^ d[8])) & (!(c[8] & d[8])) & a[7]);
    assign c[7] = ((c[8] ^ d[8]) & (! a[7]) & b[7]) | ((!(c[8] ^ d[8])) & c[8] & d[8] & 1) | ((!(c[8] ^ d[8])) & (!(c[8] & d[8])) & 0);
    assign d[7] = ((c[8] ^ d[8]) & ((! a[7]) | b[7])) | ((!(c[8] ^ d[8])) & c[8] & d[8] & 1) | ((!(c[8] ^ d[8])) & (!(c[8] & d[8])) & 0);
    
    assign answer[6] = ((c[7] ^ d[7]) & (a[6] | b[6])) | ((!(c[7] ^ d[7])) & c[7] & d[7] & b[6]) | ((!(c[7] ^ d[7])) & (!(c[7] & d[7])) & a[6]);
    assign c[6] = ((c[7] ^ d[7]) & (! a[6]) & b[6]) | ((!(c[7] ^ d[7])) & c[7] & d[7] & 1) | ((!(c[7] ^ d[7])) & (!(c[7] & d[7])) & 0);
    assign d[6] = ((c[7] ^ d[7]) & ((! a[6]) | b[6])) | ((!(c[7] ^ d[7])) & c[7] & d[7] & 1) | ((!(c[7] ^ d[7])) & (!(c[7] & d[7])) & 0);
    
    assign answer[5] = ((c[6] ^ d[6]) & (a[5] | b[5])) | ((!(c[6] ^ d[6])) & c[6] & d[6] & b[5]) | ((!(c[6] ^ d[6])) & (!(c[6] & d[6])) & a[5]);
    assign c[5] = ((c[6] ^ d[6]) & (! a[5]) & b[5]) | ((!(c[6] ^ d[6])) & c[6] & d[6] & 1) | ((!(c[6] ^ d[6])) & (!(c[6] & d[6])) & 0);
    assign d[5] = ((c[6] ^ d[6]) & ((! a[5]) | b[5])) | ((!(c[6] ^ d[6])) & c[6] & d[6] & 1) | ((!(c[6] ^ d[6])) & (!(c[6] & d[6])) & 0);
    
    assign answer[4] = ((c[5] ^ d[5]) & (a[4] | b[4])) | ((!(c[5] ^ d[5])) & c[5] & d[5] & b[4]) | ((!(c[5] ^ d[5])) & (!(c[5] & d[5])) & a[4]);
    assign c[4] = ((c[5] ^ d[5]) & (! a[4]) & b[4]) | ((!(c[5] ^ d[5])) & c[5] & d[5] & 1) | ((!(c[5] ^ d[5])) & (!(c[5] & d[5])) & 0);
    assign d[4] = ((c[5] ^ d[5]) & ((! a[4]) | b[4])) | ((!(c[5] ^ d[5])) & c[5] & d[5] & 1) | ((!(c[5] ^ d[5])) & (!(c[5] & d[5])) & 0);
    
    assign answer[3] = ((c[4] ^ d[4]) & (a[3] | b[3])) | ((!(c[4] ^ d[4])) & c[4] & d[4] & b[3]) | ((!(c[4] ^ d[4])) & (!(c[4] & d[4])) & a[3]);
    assign c[3] = ((c[4] ^ d[4]) & (! a[3]) & b[3]) | ((!(c[4] ^ d[4])) & c[4] & d[4] & 1) | ((!(c[4] ^ d[4])) & (!(c[4] & d[4])) & 0);
    assign d[3] = ((c[4] ^ d[4]) & ((! a[3]) | b[3])) | ((!(c[4] ^ d[4])) & c[4] & d[4] & 1) | ((!(c[4] ^ d[4])) & (!(c[4] & d[4])) & 0);
    
    assign answer[2] = ((c[3] ^ d[3]) & (a[2] | b[2])) | ((!(c[3] ^ d[3])) & c[3] & d[3] & b[2]) | ((!(c[3] ^ d[3])) & (!(c[3] & d[3])) & a[2]);
    assign c[2] = ((c[3] ^ d[3]) & (! a[2]) & b[2]) | ((!(c[3] ^ d[3])) & c[3] & d[3] & 1) | ((!(c[3] ^ d[3])) & (!(c[3] & d[3])) & 0);
    assign d[2] = ((c[3] ^ d[3]) & ((! a[2]) | b[2])) | ((!(c[3] ^ d[3])) & c[3] & d[3] & 1) | ((!(c[3] ^ d[3])) & (!(c[3] & d[3])) & 0);
    
    assign answer[1] = ((c[2] ^ d[2]) & (a[1] | b[1])) | ((!(c[2] ^ d[2])) & c[2] & d[2] & b[1]) | ((!(c[2] ^ d[2])) & (!(c[2] & d[2])) & a[1]);
    assign c[1] = ((c[2] ^ d[2]) & (! a[1]) & b[1]) | ((!(c[2] ^ d[2])) & c[2] & d[2] & 1) | ((!(c[2] ^ d[2])) & (!(c[2] & d[2])) & 0);
    assign d[1] = ((c[2] ^ d[2]) & ((! a[1]) | b[1])) | ((!(c[2] ^ d[2])) & c[2] & d[2] & 1) | ((!(c[2] ^ d[2])) & (!(c[2] & d[2])) & 0);
    
    assign answer[0] = ((c[1] ^ d[1]) & (a[0] | b[0])) | ((!(c[1] ^ d[1])) & c[1] & d[1] & b[0]) | ((!(c[1] ^ d[1])) & (!(c[1] & d[1])) & a[0]);
endmodule



